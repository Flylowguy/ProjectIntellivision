LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY something IS

END something;

ARCHITECTURE behaviour OF something IS
BEGIN

END behaviour;
