
LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY work;

ENTITY ALU IS
	PORT
	(
		a_inv :  IN  STD_LOGIC;
		b_inv :  IN  STD_LOGIC;
		A :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		alu_op :  IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		B :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		ZEROIN :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		C :  OUT  STD_LOGIC;
		N :  OUT  STD_LOGIC;
		V :  OUT  STD_LOGIC;
		Z :  OUT  STD_LOGIC;
		fOut :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END ALU;

ARCHITECTURE bdf_type OF ALU IS

COMPONENT rcadder
	PORT(cIn : IN STD_LOGIC;
		 aIn : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 bIn : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 c30 : OUT STD_LOGIC;
		 c31 : OUT STD_LOGIC;
		 f : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT not32
	PORT(A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 output : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mux2
	PORT(sel : IN STD_LOGIC;
		 d0 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 d1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 f : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT or32
	PORT(A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 output : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT and32
	PORT(A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 output : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT zeroflag
	PORT(A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 output : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT mux4
	PORT(d0 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 d1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 d2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 d3 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 sel : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 f : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT xor32
	PORT(A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 output : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	addAin :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	addBin :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	f :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	sel :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	zin :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC_VECTOR(31 DOWNTO 0);


BEGIN
C <= SYNTHESIZED_WIRE_2;



b2v_inst : rcadder
PORT MAP(cIn => SYNTHESIZED_WIRE_0,
		 aIn => addAin,
		 bIn => addBin,
		 c30 => SYNTHESIZED_WIRE_1,
		 c31 => SYNTHESIZED_WIRE_2,
		 f => f);


V <= SYNTHESIZED_WIRE_1 XOR SYNTHESIZED_WIRE_2;


b2v_inst11 : not32
PORT MAP(A => B,
		 output => SYNTHESIZED_WIRE_3);


b2v_inst12 : mux2
PORT MAP(sel => b_inv,
		 d0 => B,
		 d1 => SYNTHESIZED_WIRE_3,
		 f => addBin);


b2v_inst13 : or32
PORT MAP(A => addAin,
		 B => addBin,
		 output => SYNTHESIZED_WIRE_5);


b2v_inst14 : and32
PORT MAP(A => addAin,
		 B => addBin,
		 output => SYNTHESIZED_WIRE_6);


b2v_inst2 : zeroflag
PORT MAP(A => f,
		 output => Z);


SYNTHESIZED_WIRE_0 <= a_inv XOR b_inv;


b2v_inst4 : mux4
PORT MAP(d0 => f,
		 d1 => SYNTHESIZED_WIRE_4,
		 d2 => SYNTHESIZED_WIRE_5,
		 d3 => SYNTHESIZED_WIRE_6,
		 sel => sel,
		 f => fOut);


b2v_inst6 : mux2
PORT MAP(sel => a_inv,
		 d0 => A,
		 d1 => SYNTHESIZED_WIRE_7,
		 f => addAin);


b2v_inst8 : not32
PORT MAP(A => A,
		 output => SYNTHESIZED_WIRE_7);


b2v_inst9 : xor32
PORT MAP(A => addAin,
		 B => addBin,
		 output => SYNTHESIZED_WIRE_4);

N <= f(31);
sel <= alu_op;

END bdf_type;
